interface intr;
  logic I0;
  logic I1;
  logic I2;
  logic I3;
  logic a,b;
endinterface