class transaction;
  randc bit I0;
  randc bit I1;
  randc bit I2;
  randc bit I3;
  bit a,b;
endclass
